-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.0 Build 156 04/24/2013 SJ Full Version
-- Created on Mon Feb 15 20:14:59 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY project2fsm IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Key1 : IN STD_LOGIC := '0';
        Key2 : IN STD_LOGIC := '0';
        StatusA : OUT STD_LOGIC;
        StatusB : OUT STD_LOGIC
    );
END project2fsm;

ARCHITECTURE BEHAVIOR OF project2fsm IS
    TYPE type_fstate IS (Init,Test,Pause,Gen);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Key1,Key2)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Init;
            StatusA <= '0';
            StatusB <= '0';
        ELSE
            StatusA <= '0';
            StatusB <= '0';
            CASE fstate IS
                WHEN Init =>
                    reg_fstate <= Test;

                    StatusB <= '0';

                    StatusA <= '0';
                WHEN Test =>
                    IF (((Key1 = '1') AND NOT((Key2 = '1')))) THEN
                        reg_fstate <= Pause;
                    ELSIF ((NOT((Key1 = '1')) AND (Key2 = '1'))) THEN
                        reg_fstate <= Gen;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Test;
                    END IF;

                    StatusB <= '1';

                    StatusA <= '0';
                WHEN Pause =>
                    IF (((Key1 = '1') AND NOT((Key2 = '1')))) THEN
                        reg_fstate <= Test;
                    ELSIF ((NOT((Key1 = '1')) AND (Key2 = '1'))) THEN
                        reg_fstate <= Gen;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Pause;
                    END IF;

                    StatusB <= '0';

                    StatusA <= '1';
                WHEN Gen =>
                    IF ((NOT((Key1 = '1')) AND (Key2 = '1'))) THEN
                        reg_fstate <= Test;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Gen;
                    END IF;

                    StatusB <= '1';

                    StatusA <= '1';
                WHEN OTHERS => 
                    StatusA <= 'X';
                    StatusB <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
